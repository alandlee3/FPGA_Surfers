`timescale 1ns / 1ps
`default_nettype none

module tile_painter (
        input wire clk,
        input wire rst,
        input wire 
    );


endmodule

`default_nettype wire
